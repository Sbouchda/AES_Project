library ieee;
use ieee.std_logic_1164.all;

entity SubByte is
    port(
        INP  : in  std_logic_vector(7 downto 0);
        OUTP : out std_logic_vector(7 downto 0)
    );
end entity;

architecture SubByteArch of SubByte is
begin
    process(INP)
    begin
        case(INP) is
            when x"00" => OUTP <= x"63";
            when x"01" => OUTP <= x"7c";
            when x"02" => OUTP <= x"77";
            when x"03" => OUTP <= x"7b";
            when x"04" => OUTP <= x"f2";
            when x"05" => OUTP <= x"6b";
            when x"06" => OUTP <= x"6f";
            when x"07" => OUTP <= x"c5";
            when x"08" => OUTP <= x"30";
            when x"09" => OUTP <= x"01";
            when x"0a" => OUTP <= x"67";
            when x"0b" => OUTP <= x"2b";
            when x"0c" => OUTP <= x"fe";
            when x"0d" => OUTP <= x"d7";
            when x"0e" => OUTP <= x"ab";
            when x"0f" => OUTP <= x"76";
            when x"10" => OUTP <= x"ca";
            when x"11" => OUTP <= x"82";
            when x"12" => OUTP <= x"c9";
            when x"13" => OUTP <= x"7d";
            when x"14" => OUTP <= x"fa";
            when x"15" => OUTP <= x"59";
            when x"16" => OUTP <= x"47";
            when x"17" => OUTP <= x"f0";
            when x"18" => OUTP <= x"ad";
            when x"19" => OUTP <= x"d4";
            when x"1a" => OUTP <= x"a2";
            when x"1b" => OUTP <= x"af";
            when x"1c" => OUTP <= x"9c";
            when x"1d" => OUTP <= x"a4";
            when x"1e" => OUTP <= x"72";
            when x"1f" => OUTP <= x"c0";
            when x"20" => OUTP <= x"b7";
            when x"21" => OUTP <= x"fd";
            when x"22" => OUTP <= x"93";
            when x"23" => OUTP <= x"26";
            when x"24" => OUTP <= x"36";
            when x"25" => OUTP <= x"3f";
            when x"26" => OUTP <= x"f7";
            when x"27" => OUTP <= x"cc";
            when x"28" => OUTP <= x"34";
            when x"29" => OUTP <= x"a5";
            when x"2a" => OUTP <= x"e5";
            when x"2b" => OUTP <= x"f1";
            when x"2c" => OUTP <= x"71";
            when x"2d" => OUTP <= x"d8";
            when x"2e" => OUTP <= x"31";
            when x"2f" => OUTP <= x"15";
            when x"30" => OUTP <= x"04";
            when x"31" => OUTP <= x"c7";
            when x"32" => OUTP <= x"23";
            when x"33" => OUTP <= x"c3";
            when x"34" => OUTP <= x"18";
            when x"35" => OUTP <= x"96";
            when x"36" => OUTP <= x"05";
            when x"37" => OUTP <= x"9a";
            when x"38" => OUTP <= x"07";
            when x"39" => OUTP <= x"12";
            when x"3a" => OUTP <= x"80";
            when x"3b" => OUTP <= x"e2";
            when x"3c" => OUTP <= x"eb";
            when x"3d" => OUTP <= x"27";
            when x"3e" => OUTP <= x"b2";
            when x"3f" => OUTP <= x"75";
            when x"40" => OUTP <= x"09";
            when x"41" => OUTP <= x"83";
            when x"42" => OUTP <= x"2c";
            when x"43" => OUTP <= x"1a";
            when x"44" => OUTP <= x"1b";
            when x"45" => OUTP <= x"6e";
            when x"46" => OUTP <= x"5a";
            when x"47" => OUTP <= x"a0";
            when x"48" => OUTP <= x"52";
            when x"49" => OUTP <= x"3b";
            when x"4a" => OUTP <= x"d6";
            when x"4b" => OUTP <= x"b3";
            when x"4c" => OUTP <= x"29";
            when x"4d" => OUTP <= x"e3";
            when x"4e" => OUTP <= x"2f";
            when x"4f" => OUTP <= x"84";
            when x"50" => OUTP <= x"53";
            when x"51" => OUTP <= x"d1";
            when x"52" => OUTP <= x"00";
            when x"53" => OUTP <= x"ed";
            when x"54" => OUTP <= x"20";
            when x"55" => OUTP <= x"fc";
            when x"56" => OUTP <= x"b1";
            when x"57" => OUTP <= x"5b";
            when x"58" => OUTP <= x"6a";
            when x"59" => OUTP <= x"cb";
            when x"5a" => OUTP <= x"be";
            when x"5b" => OUTP <= x"39";
            when x"5c" => OUTP <= x"4a";
            when x"5d" => OUTP <= x"4c";
            when x"5e" => OUTP <= x"58";
            when x"5f" => OUTP <= x"cf";
            when x"60" => OUTP <= x"d0";
            when x"61" => OUTP <= x"ef";
            when x"62" => OUTP <= x"aa";
            when x"63" => OUTP <= x"fb";
            when x"64" => OUTP <= x"43";
            when x"65" => OUTP <= x"4d";
            when x"66" => OUTP <= x"33";
            when x"67" => OUTP <= x"85";
            when x"68" => OUTP <= x"45";
            when x"69" => OUTP <= x"f9";
            when x"6a" => OUTP <= x"02";
            when x"6b" => OUTP <= x"7f";
            when x"6c" => OUTP <= x"50";
            when x"6d" => OUTP <= x"3c";
            when x"6e" => OUTP <= x"9f";
            when x"6f" => OUTP <= x"a8";
            when x"70" => OUTP <= x"51";
            when x"71" => OUTP <= x"a3";
            when x"72" => OUTP <= x"40";
            when x"73" => OUTP <= x"8f";
            when x"74" => OUTP <= x"92";
            when x"75" => OUTP <= x"9d";
            when x"76" => OUTP <= x"38";
            when x"77" => OUTP <= x"f5";
            when x"78" => OUTP <= x"bc";
            when x"79" => OUTP <= x"b6";
            when x"7a" => OUTP <= x"da";
            when x"7b" => OUTP <= x"21";
            when x"7c" => OUTP <= x"10";
            when x"7d" => OUTP <= x"ff";
            when x"7e" => OUTP <= x"f3";
            when x"7f" => OUTP <= x"d2";
            when x"80" => OUTP <= x"cd";
            when x"81" => OUTP <= x"0c";
            when x"82" => OUTP <= x"13";
            when x"83" => OUTP <= x"ec";
            when x"84" => OUTP <= x"5f";
            when x"85" => OUTP <= x"97";
            when x"86" => OUTP <= x"44";
            when x"87" => OUTP <= x"17";
            when x"88" => OUTP <= x"c4";
            when x"89" => OUTP <= x"a7";
            when x"8a" => OUTP <= x"7e";
            when x"8b" => OUTP <= x"3d";
            when x"8c" => OUTP <= x"64";
            when x"8d" => OUTP <= x"5d";
            when x"8e" => OUTP <= x"19";
            when x"8f" => OUTP <= x"73";
            when x"90" => OUTP <= x"60";
            when x"91" => OUTP <= x"81";
            when x"92" => OUTP <= x"4f";
            when x"93" => OUTP <= x"dc";
            when x"94" => OUTP <= x"22";
            when x"95" => OUTP <= x"2a";
            when x"96" => OUTP <= x"90";
            when x"97" => OUTP <= x"88";
            when x"98" => OUTP <= x"46";
            when x"99" => OUTP <= x"ee";
            when x"9a" => OUTP <= x"b8";
            when x"9b" => OUTP <= x"14";
            when x"9c" => OUTP <= x"de";
            when x"9d" => OUTP <= x"5e";
            when x"9e" => OUTP <= x"0b";
            when x"9f" => OUTP <= x"db";
            when x"a0" => OUTP <= x"e0";
            when x"a1" => OUTP <= x"32";
            when x"a2" => OUTP <= x"3a";
            when x"a3" => OUTP <= x"0a";
            when x"a4" => OUTP <= x"49";
            when x"a5" => OUTP <= x"06";
            when x"a6" => OUTP <= x"24";
            when x"a7" => OUTP <= x"5c";
            when x"a8" => OUTP <= x"c2";
            when x"a9" => OUTP <= x"d3";
            when x"aa" => OUTP <= x"ac";
            when x"ab" => OUTP <= x"62";
            when x"ac" => OUTP <= x"91";
            when x"ad" => OUTP <= x"95";
            when x"ae" => OUTP <= x"e4";
            when x"af" => OUTP <= x"79";
            when x"b0" => OUTP <= x"e7";
            when x"b1" => OUTP <= x"c8";
            when x"b2" => OUTP <= x"37";
            when x"b3" => OUTP <= x"6d";
            when x"b4" => OUTP <= x"8d";
            when x"b5" => OUTP <= x"d5";
            when x"b6" => OUTP <= x"4e";
            when x"b7" => OUTP <= x"a9";
            when x"b8" => OUTP <= x"6c";
            when x"b9" => OUTP <= x"56";
            when x"ba" => OUTP <= x"f4";
            when x"bb" => OUTP <= x"ea";
            when x"bc" => OUTP <= x"65";
            when x"bd" => OUTP <= x"7a";
            when x"be" => OUTP <= x"ae";
            when x"bf" => OUTP <= x"08";
            when x"c0" => OUTP <= x"ba";
            when x"c1" => OUTP <= x"78";
            when x"c2" => OUTP <= x"25";
            when x"c3" => OUTP <= x"2e";
            when x"c4" => OUTP <= x"1c";
            when x"c5" => OUTP <= x"a6";
            when x"c6" => OUTP <= x"b4";
            when x"c7" => OUTP <= x"c6";
            when x"c8" => OUTP <= x"e8";
            when x"c9" => OUTP <= x"dd";
            when x"ca" => OUTP <= x"74";
            when x"cb" => OUTP <= x"1f";
            when x"cc" => OUTP <= x"4b";
            when x"cd" => OUTP <= x"bd";
            when x"ce" => OUTP <= x"8b";
            when x"cf" => OUTP <= x"8a";
            when x"d0" => OUTP <= x"70";
            when x"d1" => OUTP <= x"3e";
            when x"d2" => OUTP <= x"b5";
            when x"d3" => OUTP <= x"66";
            when x"d4" => OUTP <= x"48";
            when x"d5" => OUTP <= x"03";
            when x"d6" => OUTP <= x"f6";
            when x"d7" => OUTP <= x"0e";
            when x"d8" => OUTP <= x"61";
            when x"d9" => OUTP <= x"35";
            when x"da" => OUTP <= x"57";
            when x"db" => OUTP <= x"b9";
            when x"dc" => OUTP <= x"86";
            when x"dd" => OUTP <= x"c1";
            when x"de" => OUTP <= x"1d";
            when x"df" => OUTP <= x"9e";
            when x"e0" => OUTP <= x"e1";
            when x"e1" => OUTP <= x"f8";
            when x"e2" => OUTP <= x"98";
            when x"e3" => OUTP <= x"11";
            when x"e4" => OUTP <= x"69";
            when x"e5" => OUTP <= x"d9";
            when x"e6" => OUTP <= x"8e";
            when x"e7" => OUTP <= x"94";
            when x"e8" => OUTP <= x"9b";
            when x"e9" => OUTP <= x"1e";
            when x"ea" => OUTP <= x"87";
            when x"eb" => OUTP <= x"e9";
            when x"ec" => OUTP <= x"ce";
            when x"ed" => OUTP <= x"55";
            when x"ee" => OUTP <= x"28";
            when x"ef" => OUTP <= x"df";
            when x"f0" => OUTP <= x"8c";
            when x"f1" => OUTP <= x"a1";
            when x"f2" => OUTP <= x"89";
            when x"f3" => OUTP <= x"0d";
            when x"f4" => OUTP <= x"bf";
            when x"f5" => OUTP <= x"e6";
            when x"f6" => OUTP <= x"42";
            when x"f7" => OUTP <= x"68";
            when x"f8" => OUTP <= x"41";
            when x"f9" => OUTP <= x"99";
            when x"fa" => OUTP <= x"2d";
            when x"fb" => OUTP <= x"0f";
            when x"fc" => OUTP <= x"b0";
            when x"fd" => OUTP <= x"54";
            when x"fe" => OUTP <= x"bb";
            when x"ff" => OUTP <= x"16";
            when others => OUTP <= (others => '0');
        end case;
    end process;
end architecture;
